
module _and_gate #(BITS=8) (
  input logic [BITS-1:0] a,
  input logic [BITS-1:0] b,
  output logic [BITS-1:0] c
);
endmodule


