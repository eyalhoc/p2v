module hello_world ();


endmodule
