module params__bits8_namefoo_sampleFalse ();

    // params module parameters:
    //  * clk = clk_arst() (p2v_clock) #  p2v clock
    //  * bits = 8 (int) #  integer parameter
    //  * name = "foo" (str) #  string parameter
    //  * sample = False (bool) #  bool parameter - no constraint
    //  * d = {} (dict) #  dictionary parameter - complex parameter does not create suffix automatcically
    //  * depth = 128 (int) #  integer parameter - does not affect module name


endmodule  // params__bits8_namefoo_sampleFalse
