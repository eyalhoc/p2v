module params__bits8_namefoo_sampleFalse ();

    // module parameters:
    // clk = p2v_clock.clk_arst() (p2v_clock)
    // bits = 8 (int)
    // name = "foo" (str)
    // sample = False (bool)
    // d = {} (dict)
    // depth = 128 (int)


endmodule
