module hello_world ();

    // hello_world module parameters:


endmodule  // hello_world
